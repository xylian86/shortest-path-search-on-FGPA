module ADD_SUB9