module  usbmouse (input         Clk,                // 50 MHz clock
                             Reset,              // Active-high reset signal
                             frame_clk,          // The clock indicating a new frame (~60Hz)
               input [9:0]   DrawX, DrawY,       // Current pixel coordinates
					input logic [7:0] keycode,
					input logic STOREBEGIN,STOREEND,
               output logic  is_ball,is_usbmouse,          // Whether current pixel belongs to ball or background
					output logic [9:0] Ball_X_OUT, Ball_Y_OUT
              );
    
    parameter [9:0] Ball_X_Center = 10'd320;  // Center position on the X axis
    parameter [9:0] Ball_Y_Center = 10'd240;  // Center position on the Y axis
    parameter [9:0] Ball_X_Min = 10'd0;       // Leftmost point on the X axis
    parameter [9:0] Ball_X_Max = 10'd639;     // Rightmost point on the X axis
    parameter [9:0] Ball_Y_Min = 10'd0;       // Topmost point on the Y axis
    parameter [9:0] Ball_Y_Max = 10'd479;     // Bottommost point on the Y axis
    parameter [9:0] Ball_X_Step = 10'd1;      // Step size on the X axis
    parameter [9:0] Ball_Y_Step = 10'd1;      // Step size on the Y axis
    parameter [9:0] Ball_Size = 10'd3;        // Ball size
    
    logic [9:0] Ball_X_Pos, Ball_X_Motion, Ball_Y_Pos, Ball_Y_Motion;
    logic [9:0] Ball_X_Pos_in, Ball_X_Motion_in, Ball_Y_Pos_in, Ball_Y_Motion_in;
	 logic [7:0] w,a,s,d,space;
	 
	 logic [9:0] BEGINX,BEGINY,ENDX,ENDY;
	 
	 assign w=8'b00011010;
	 assign a=8'b00000100;
	 assign s=8'b00010110;
	 assign d=8'b00000111;
	 assign space=8'h2c;
	 
	 assign Ball_X_OUT=Ball_X_Pos;
	 assign Ball_Y_OUT=Ball_Y_Pos;
    
    //////// Do not modify the always_ff blocks. ////////
    // Detect rising edge of frame_clk
    logic frame_clk_delayed, frame_clk_rising_edge;
    always_ff @ (posedge Clk) begin
        frame_clk_delayed <= frame_clk;
        frame_clk_rising_edge <= (frame_clk == 1'b1) && (frame_clk_delayed == 1'b0);
    end
    // Update registers
	 always_ff @ (STOREBEGIN)
	 begin
	 BEGINX<=Ball_X_Pos;
	 BEGINY<=Ball_Y_Pos;
	 end
	 
	 always_ff @ (STOREEND)
	 begin
	 ENDX<=Ball_X_Pos;
	 ENDY<=Ball_Y_Pos;
	 end
	  
    always_ff @ (posedge Clk)
    begin
        if (Reset)
        begin
            Ball_X_Pos <= Ball_X_Center;
            Ball_Y_Pos <= Ball_Y_Center;
            Ball_X_Motion <= 10'd0;
            Ball_Y_Motion <= 10'd0;
        end
        else
        begin
            Ball_X_Pos <= Ball_X_Pos_in;
            Ball_Y_Pos <= Ball_Y_Pos_in;
            Ball_X_Motion <= Ball_X_Motion_in;
            Ball_Y_Motion <= Ball_Y_Motion_in;
        end
    end
    //////// Do not modify the always_ff blocks. ////////
    
    // You need to modify always_comb block.
    always_comb
    begin
        // By default, keep Motion and position unchanged
        Ball_X_Pos_in = Ball_X_Pos;
        Ball_Y_Pos_in = Ball_Y_Pos;
        Ball_X_Motion_in = Ball_X_Motion;
        Ball_Y_Motion_in = Ball_Y_Motion;
        
        // Update position and Motion only at rising edge of frame clock
        if (frame_clk_rising_edge)
        begin
            // Be careful when using comparators with "logic" datatype because compiler treats 
            //   both sides of the operator as UNSIGNED numbers.
            // e.g. Ball_Y_Pos - Ball_Size <= Ball_Y_Min 
            // If Ball_Y_Pos is 0, then Ball_Y_Pos - Ball_Size will not be -4, but rather a large positive number.
            // Pay attention to the velocity. We must always make sure that the ball only has velocity in one direction.
				if (keycode==w)
					begin
						Ball_Y_Motion_in=(~(Ball_Y_Step)+1'b1);
						Ball_X_Motion_in=10'd0;
					end
				else if (keycode==a)
					begin
						Ball_X_Motion_in=(~(Ball_X_Step)+1'b1);
						Ball_Y_Motion_in=10'd0;
					end
				else if (keycode==s)
					begin
						Ball_Y_Motion_in=Ball_Y_Step;
						Ball_X_Motion_in=10'd0;
					end
				else if (keycode==d)
					begin
						Ball_X_Motion_in=Ball_X_Step;
						Ball_Y_Motion_in=10'd0;
					end
				else if (keycode==8'd0)
					begin
						Ball_X_Motion_in=10'd0;
						Ball_Y_Motion_in=10'd0;
					end
				
			
//				//Update part
//				if( Ball_Y_Pos + Ball_Size >= Ball_Y_Max )  // Ball is at the bottom edge, BOUNCE!
//					begin
//						Ball_Y_Motion_in = (~(Ball_Y_Step) + 1'b1);  // 2's complement.  
//						Ball_X_Motion_in=10'd0;
//					end
//            else if ( Ball_Y_Pos <= Ball_Y_Min + Ball_Size )  // Ball is at the top edge, BOUNCE!
//                begin
//						Ball_Y_Motion_in = Ball_Y_Step;
//						Ball_X_Motion_in=10'd0;
//					 end
//            // TODO: Add other boundary detections and handle keypress here.
//				else if( Ball_X_Pos + Ball_Size >= Ball_X_Max )  // Ball is at the right edge, BOUNCE!
//					begin
//						Ball_X_Motion_in = (~(Ball_X_Step) + 1'b1);  // 2's complement.  
//						Ball_Y_Motion_in=10'd0;
//					end
//            else if ( Ball_X_Pos <= Ball_X_Min + Ball_Size )  // Ball is at the left edge, BOUNCE!
//                begin
//						Ball_X_Motion_in = Ball_X_Step;
//						Ball_Y_Motion_in=10'd0;
//					 end
        
            // Update the ball's position with its Motion
            Ball_X_Pos_in = Ball_X_Pos + Ball_X_Motion;
            Ball_Y_Pos_in = Ball_Y_Pos + Ball_Y_Motion;
        end
        
        /**************************************************************************************
            ATTENTION! Please answer the following quesiton in your lab report! Points will be allocated for the answers!
            Hidden Question #2/2:
               Notice that Ball_Y_Pos is updated using Ball_Y_Motion. 
              Will the new value of Ball_Y_Motion be used when Ball_Y_Pos is updated, or the old? 
              What is the difference between writing
                "Ball_Y_Pos_in = Ball_Y_Pos + Ball_Y_Motion;" and 
                "Ball_Y_Pos_in = Ball_Y_Pos + Ball_Y_Motion_in;"?
              How will this impact behavior of the ball during a bounce, and how might that interact with a response to a keypress?
              Give an answer in your Post-Lab.
				Answer:1. It has been updated when Ball_Y_Pos is updated. 2. For the design "Ball_Y_Pos_in = Ball_Y_Pos + Ball_Y_Motion;" ,
				The frame will create one delay so that the ball will go through the boundary for a while and then back to the screen; for the design "Ball_Y_Pos_in = Ball_Y_Pos + Ball_Y_Motion_in;",
				The ball will response the keyboard immediately and there will be no frame delay for the ball moving.
        **************************************************************************************/
    end
    
    // Compute whether the pixel corresponds to ball or background
    /* Since the multiplicants are required to be signed, we have to first cast them
       from logic to int (signed by default) before they are multiplied. */
    int DistX, DistY, Size;
    assign DistX = DrawX - Ball_X_Pos;
    assign DistY = DrawY - Ball_Y_Pos;
    assign Size = Ball_Size;
    always_comb begin
        if ( ( DistX*DistX + DistY*DistY) <= (Size*Size) ) 
            is_usbmouse = 1'b1;
        else
            is_usbmouse = 1'b0;
        /* The ball's (pixelated) circle is generated using the standard circle formula.  Note that while 
           the single line is quite powerful descriptively, it causes the synthesis tool to use up three
           of the 12 available multipliers on the chip! */
    end
    
endmodule