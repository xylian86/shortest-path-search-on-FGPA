module ramstore4(input [9:0] DrawX, DrawY, output [1:0] data4);       // Current pixel coordinates

//begin graph
parameter [479:0][639:0][1:0] maplist={{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,},
{2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,},
{2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,},
{2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,},
{2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,},
{2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,},
{2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,},
{2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,},
{2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,},
{2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,},
{2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,},
{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,},
{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,},
{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,},
{2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,},
{2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,},
{2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,},
{2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,},
{2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,},
{2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,},
{2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,},
{2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,},
{2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,},
{2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,},
{2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,},
{2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,},
{2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,},
{2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,},
{2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd2,2'd0,},
{2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,},
{2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,},
{2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,},
{2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd1,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd1,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,},
{2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,},
{2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd1,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd1,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd1,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd1,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd1,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,},
{2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd1,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd2,2'd0,2'd0,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd1,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,},
{2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,},
{2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,},
{2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,},
{2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,},
{2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,},
{2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,},
{2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,},
{2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,},
{2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,},
{2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,},
{2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,},
{2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,},
{2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,},
{2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,},
{2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,},
{2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,},
{2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,},
{2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,},
{2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd1,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,},
{2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,},
{2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,},
{2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,},
{2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,},
{2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,},
{2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,},
{2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd1,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,},
{2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,},
{2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,},
{2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,},
{2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,},
{2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd1,2'd0,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd1,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,},
{2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,},
{2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd1,2'd2,2'd0,2'd1,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,},
{2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,},
{2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd2,2'd2,2'd1,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,},
{2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd1,2'd1,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,},
{2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd2,2'd1,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,},
{2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd1,2'd2,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,},
{2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd1,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,},
{2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,},
{2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,},
{2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,},
{2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,},
{2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,},
{2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,},
{2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd1,2'd1,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,},
{2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,},
{2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd0,2'd0,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,},
{2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd1,2'd1,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,},
{2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd0,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd1,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd2,2'd1,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd1,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd1,2'd2,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd2,2'd0,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,},
{2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,},
{2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd1,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,},
{2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd0,2'd2,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,},
{2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd2,2'd0,2'd2,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,},
{2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,},
{2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},
{2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,},};


always_comb
	begin
		if (DrawX<10'd640 && DrawY<10'd480)
		begin
			data4=maplist[10'd479-DrawY][10'd639-DrawX];
		end
		else
		begin
			data4=2'd0;
		end
	end
endmodule